module Example03_using_wand(a,b,c,d,f);
  input a,b,c,d;
  output wand f;
  assign f = a&b;
  assign f = c|d;
endmodule 
