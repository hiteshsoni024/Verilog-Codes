module Example03_using_wor(a,b,c,d,f);
  input a,b,c,d;
  output wor f;
  assign f = a&b;
  assign f = c|d;
endmodule 
